// note the original should contain 4 buffers = 2 in, 2 out = each of 512 bytes (it corresponds to fpga_flash_fifo in versatile_fifo docs)
// then we also try to make only 2 buffers - one in, one out
// original prefixes were w b _ (Wishbone) and s d _ (SD card)
// then we rename to u s b f t _ (FTDI USB) and f p g a _ (FPGA internal) , respectively...
// NOW, here we have but one buffer - writable from one side, readable from other, with different clock domains.
// so instead of u s b f t _ and f p g a _ , will refer to r d _ and w r _ sides of the buffer..

module versatile_sd_fifo_1buf
  (
    input [7:0]  dat_i, // data input
    output [7:0] dat_o, // data output
    input 	 we_i, // write enable input - works only on wr_clk
    input 	 re_i, //read enable input -  works only on rd_clk
    input 	 wr_clk,
    input 	 rd_clk, // one buffer, but we leave this since we want dual clock

    output fifo_full, // only one buffer
    output fifo_empty, // only one buffer
    output fifo_aempty, // only one buffer - "asynchron" empty (quicker)
    input 	 rst
  );


  //buffering the clocks - to clear out (*) These 2 clock signal(s) are generated by combinatorial logic ... ambiguities?
  // wire w_clk, r_clk;
  // wire wr_clk_buf, rd_clk_buf;

  // IBUFG r_buf_1 ( .O(rd_clk_buf), .I (rd_clk) );
  // BUFG r_buf_2 ( .O (r_clk), .I (rd_clk_buf) );//For best clock quality

  // IBUFG w_buf_1 ( .O(wr_clk_buf), .I (wr_clk) );
  // BUFG w_buf_2 ( .O (w_clk), .I (wr_clk_buf) );//For best clock quality


  // only one buffer now - but keep the "1" suffixes
  // orig 9 bit - [8:0] for .ADDR_WIDTH(9)
  wire [8:0] 	 wptr1, rptr1; // write, read pointer
  wire [8:0] 	 wadr1, radr1; // write, read address

  wire 	 dpram_we_a;
  //wire [9:0] 	 dpram_a_a, dpram_a_b;   // dpram address wire [9:0] for  .ADDR_WIDTH(9) - only one buffer now, not 10 bit wide (no address selector)
  wire [8:0] 	 dpram_a_a;   // dpram address - only one buffer now, but these are write & read addresses //9 bit
  wire [8:0] 	 dpram_a_b;
  wire [7:0] 	 wdat_o; // seems need to define wire for a proper connection to RAM out

  wire rstplus;
  reg rstplusR; //was wire - do not init these
  reg rstplusR2;

  // replacement variables for cke contructs below
  wire wptr_en;
  wire rptr_en;
  reg wptr_en_once; //'one-shot'-ted; cannot be wire if set in FSM
  reg wonce_state;
  reg rptr_en_once; //'one-shot'-ted; cannot be wire if set in FSM
  reg ronce_state;

  initial begin
    wonce_state=0;
    ronce_state=0;
    // "Reference to vector wire 'wadr1' is not a legal reg or variable lvalue"
    // fixed init by changing CNT_RESET_VALUE in versatile_sd_counter;
    // wptr1 = 9'b0; rptr1 = 9'b0; wadr1 = 9'b0; radr1 = 9'b0;
  end

  // mind the mixup here: if we get re_i, there is byte to read from FT,
  //   which means we want to write it to our RAM,
  //   unless the fifo is *full*!
  // Hence, do *not* use rptr_en=(re_i & !fifo_aempty); - use full there!
  // same for wptr!
	assign rptr_en = (re_i & !fifo_full);
	assign wptr_en = (we_i & !fifo_aempty);

  // eeh... note: 'dpram_we_a' IS 'rptr_en'; and 'dpram_re_b' IS 'wptr_en'
  // wire we_i = 1'bz; // repeat for port - 'Illegal redeclaration'
  //~ reg we_i = 1'bz; // repeat for port - 'Illegal redeclaration'
  // again - if this write enable - use not empty (not "(!fifo_full)" !!)
	assign dpram_we_a = (!fifo_aempty) ? we_i : 1'b0; // this gets automatically compacted with .cke(we_i & !fifo_full),
	assign dpram_a_a = wadr1; //strictly write address

   // only one buffer now - but still need this - read address
	assign dpram_a_b = radr1;
	//assign dpram_re_b = (!fifo_empty) ? re_i : 1'b0; // added - should get automatically compacted with .cke(re_i & !fifo_empty)

	//assign rstplus = (rst || fifo_full);
	//assign rstplus = (!fifo_full) ? rst : 1'b1; // here rstplus is wire; cannot do "(!fifo_full) ? 1'b0 : 1'b1;" cuz we need rst too - so seems it must be clocked
	assign rstplus = (rst || rstplusR);

  // need this continuous assignment too - else wire and port are not connected!
  assign dat_o = wdat_o;

  versatile_sd_counter wptr1_cnt
  (
    .q(wptr1),		// goes to async cmp
    .q_bin(wadr1), // dpram_a_a =wadr1;
    .cke(wptr_en_once), // was wptr_en
    .clk(wr_clk), // was wr_clk
    .rst(rstplus)
  );

  versatile_sd_counter rptr1_cnt
  (
    .q(rptr1),
    .q_bin(radr1),
    .cke(rptr_en_once), // was rptr_en; was .cke(re_i & !fifo_empty),
    .clk(rd_clk), //was rd_clk
    .rst(rstplus)
  );

  versatile_fifo_async_cmp
  #
  (
    .ADDR_WIDTH(9) //was for two buffers 9
  )
  cmp1
  (
    //.wptr(wptr1),
    .wptr(wadr1),
    //.rptr(rptr1),
    .rptr(radr1),
    .fifo_empty(fifo_empty),
    .fifo_aempty(fifo_aempty),
    .fifo_full(fifo_full),
    .wclk(wr_clk), // was wr_clk
    .rclk(rd_clk), // was rd_clk
    .rst(rstplus)
  );

   //only one buffer now - but still want it dual clock.. - so use vfifo_dual_port_ram_dc_sw
  vfifo_dual_port_ram_dc_sw
  #
  (
    // .ADDR_WIDTH(10), //only one buffer now, no concatenation in  assign dpram_a_ - address goes direct
    .ADDR_WIDTH(9),
    .DATA_WIDTH(8)
  )/* */
  dpram
  (
    .d_a(dat_i), // strictly write data in
    .adr_a(dpram_a_b),  //strictly write address - dpram_a_a=wadr1
                        // but as we're clocked with rptr now;
                        // use dpram_a_b=radr1 which changes with that clock
    .we_a(rptr_en), // write enable - only on (posedge clk_a);
                    // was: dpram_we_a - but we write to RAM,
                    //  when there is something to read from FT245!
    .clk_a(wr_clk),  // "write" clock, was usbft_clk, was wr_clk
    .q_b(wdat_o), // strictly read data out
    .adr_b(dpram_a_a), // strictly read address  - dpram_a_b=radr1
                        // but as we're clocked with wptr now;
                        // use dpram_a_a=wadr1 which changes with that clock
    //.re_b(dpram_we_b), // read enable - only on (posedge clk_b) // added bonus to prevent XX reads..
    // going back to read enable - to ensure proper transitions?
    .re_b(wptr_en), // we read from RAM only when FPGA wants to write to FT245!
    .clk_b(rd_clk) // "read" clock, was fpga_clk, was rd_clk
  );

  // 'one-shot' state machines
  // - to avoid multiple clocking of indexes, when
  // - signals come in for read & write
  always @ (posedge wr_clk)
  begin: fsm_wonce
    case (wonce_state)
    0 : begin
        wptr_en_once <= 0;
        if ( wptr_en == 1 )
          begin
            wonce_state <= 1;
            wptr_en_once <= 1;
          end
        else
          wonce_state <= 0;
      end

    1 : begin
        if ( wptr_en == 1 )
          begin
            wptr_en_once <= 0;
            wonce_state <= 1;
          end
        else
          wonce_state <= 2;
      end

    2: begin
        wonce_state <= 0;
        wptr_en_once <= 0;
      end
    endcase
  end

  always @ (posedge rd_clk)
  begin: fsm_ronce
    case (ronce_state)
    0 : begin
        rptr_en_once <= 0;
        if ( rptr_en == 1 )
          begin
            ronce_state <= 1;
            rptr_en_once <= 1;
          end
        else
          ronce_state <= 0;
      end

    1 : begin
        if ( rptr_en == 1 )
          begin
            rptr_en_once <= 0;
            ronce_state <= 1;
          end
        else
          ronce_state <= 2;
      end

    2: begin
        ronce_state <= 0;
        rptr_en_once <= 0;
      end
    endcase
  end

// clocked rstplus - needs to be a reg.
// wr_clk is currently gCLK for both instances, but the reading one isnt !!
// always @ (posedge wr_clk)
// begin : rstpl_clocked
// if (rst == 1'b1)
	// begin
		// rstplusR <= 1'b1; //reset when rst
	// end
// else   // rst is zero
	// begin
		// //rstplusR <= (!fifo_full) ? 1'b0 : 1'b1; //? rst : 1'b1;
		// if (fifo_full == 1'b0)
			// begin
				// rstplusR <= 1'b0 ;
			// end
		// else
			// begin
				// rstplusR <= 1'b1 ;
			// end
	// end
// end

// this doesn't seem to change the rstplus at all - but post-route streams..
always @ (posedge wr_clk or posedge rst or posedge fifo_full)
 if (rst)
   {rstplusR, rstplusR2} <= 2'b00;
 else if (fifo_full)
   {rstplusR, rstplusR2} <= 2'b11;
 else
   {rstplusR, rstplusR2} <= {rstplusR2, fifo_full};



endmodule // versatile_sd_fifo_1buf
